library IEEE;
use ieee.std_logic_1164.all;


entity multiplexador2x1 is 
   generic(largura: natural := 8);
   port(
      entrada0, entrada1: in std_logic_vector(largura-1 downto 0);
      selecao: in std_logic;
      saida: out std_logic_vector(largura-1 downto 0)
   );
end entity;

architecture comportamental of multiplexador2x1 is
begin
	saida <= entrada0 when selecao='0' else
			entrada1;
end architecture;
